work.Reg(Behavior) :32:
