cad_lib.Mux2(Behavior) :32:
cad_lib.Reg(Behavior) :32:
cad_lib.ALU(behavior) rtlc_no_parameters
cad_lib.Reg(Behavior) :5:
cad_lib.Fun_reg(Behavior) rtlc_no_parameters
cad_lib.Reg_dec(Behavior) rtlc_no_parameters
cad_lib.Mux32(Behavior) rtlc_no_parameters
