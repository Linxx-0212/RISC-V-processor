work.Mux2(Behavior) :32:
