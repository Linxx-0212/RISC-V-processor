cad_lib.Reg_dec(Behavior) rtlc_no_parameters
cad_lib.Reg(Behavior) :32:
cad_lib.Mux32(Behavior) rtlc_no_parameters
