work.Reg_dec(Behavior) rtlc_no_parameters
work.Reg(Behavior) :32:
