cad_lib.Mux2(Behavior) :32:
