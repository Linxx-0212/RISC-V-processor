work.Reg_dec(Behavior) rtlc_no_parameters
work.Reg(Behavior) :32:
work.Mux32(Behavior) rtlc_no_parameters
