work.Reg(Behavior) :32:
work.Mux2(Behavior) :32:
