work.Mux2(Behavior) :32:
work.Reg(Behavior) :32:
work.ALU(behavior) rtlc_no_parameters
work.Reg(Behavior) :5:
work.Fun_reg(Behavior) rtlc_no_parameters
work.Reg_dec(Behavior) rtlc_no_parameters
work.Mux32(Behavior) rtlc_no_parameters
