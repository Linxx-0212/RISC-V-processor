cad_lib.Reg(Behavior) :32:
